`ifndef AXI4LITEMASTERAGENT_INCLUDED_
`define AXI4LITEMASTERAGENT_INCLUDED_

module Axi4LiteMasterAgent();


endmodule: Axi4LiteMasterAgent

