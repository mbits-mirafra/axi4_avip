`ifndef AXI4LITESLAVEAGENT_INCLUDED_
`define AXI4LITESLAVEAGENT_INCLUDED_

module Axi4LiteSlaveAgent();


endmodule: Axi4LiteSlaveAgent

